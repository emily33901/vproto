module compiler

fn to_v_field_name(name string) string {
	return name.to_lower()
}

fn to_v_struct_name(name string) string {
	mut new_name := name[0].str().to_upper() + name[1..]
	new_name = new_name.replace_each(['_', '', '.', ''])

	// Get around the capital letters limitations
	mut was_cap := 0
	for i, c in new_name {
		if c >= `A` && c <= `Z` {
			if was_cap > 1 {
				new_name = new_name[..i] + c.str().to_lower() + new_name[i+1..]
			} else {
				was_cap++
			}
		} else {
			was_cap = 0
		}
	}

	return new_name
}

fn to_v_interface_name(context []string, name string) string {
	mut struct_name := ''
	
	for _, part in context {
		struct_name += to_v_struct_name(part)
	}

	struct_name += to_v_struct_name(name)

	// TODO when this limitation is removed also do so here!

	struct_name = struct_name.replace_each(['.', ''])

	return struct_name + 'er'
}

fn to_v_internal_struct_name(context []string, name string) string {
	mut struct_name := 'Internal'
	for _, part in context {
		struct_name += to_v_struct_name(part)
	}
	
	return struct_name + to_v_struct_name(name)
}

fn escape_name(name string) string {
	if name in keywords_v {
		return name + '_'
	}

	new_name := name.replace_each(['__', '_'])

	return new_name
}

struct Gen {
	type_table &TypeTable
}

fn (g &Gen) gen_file_header(f &File) string {
	// TODO figure out an appropriate module
	// if the file doesnt have an explicit package set

	return '
// Generated by vproto - Do not modify
module vproto_gen

import vproto
'
}

fn  (g &Gen) gen_enum_definition(type_context []string, e &Enum) string {
	e_name := to_v_struct_name(type_context.join('') + e.name)
	mut text := '\nenum ${e_name} {\n'

	for _, field in e.fields {
		text += '\t${to_v_field_name(field.name)} = $field.value.value\n'
	}

	text += '}\n'
	
	// TODO helper functions here 
	// https://developers.google.com/protocol-buffers/docs/reference/cpp-generated#enum

	return text
}

fn (g &Gen) type_to_type(t string, use_interface bool) (string, bool) {
	if t in valid_types {
		return valid_types_v[valid_types.index(t)], false
	}

	name_transform := if use_interface {
		to_v_interface_name
	} else {
		to_v_internal_struct_name
	}

	if _ := g.type_table.lookup_message([], t) {
		if t[0] == `.` {
			return name_transform([], t[1..]), true
		}

		return name_transform([], t), true
	}

	if t[0] == `.` {
		return to_v_struct_name(t[1..]), false
	}

	return to_v_struct_name(t), false
}

fn (g &Gen) field_type_to_type(f &Field, use_interface bool) (string, bool) {
	return g.type_to_type(f.t, use_interface)
}

fn (g &Gen) gen_message_definition(type_context []string, m &Message) string {
	mut text := ''

	m_name := to_v_interface_name(type_context, m.name)

	// Generate for submessages and subenums
	for _, e in m.enums {
		mut context := type_context
		context << m.name
		text += g.gen_enum_definition(context, e)
	}

	for _, sub in m.messages {
		mut context := type_context
		context << m.name
		text += g.gen_message_definition(context, sub)
	}


	text += '\ninterface ${m_name} { \n'

	for _, field in m.fields {
		field_type, _ := g.field_type_to_type(&field, true)
		name := escape_name(field.name)

		// TODO cleanup this whackyness when string interpolation
		// is less buggy
		
		if field.label == 'optional' || field.label == 'required' {
			text += '\t${name}() ?$field_type\n'
			text += '\tmutable_${name}() ?&$field_type\n'
			text += '\tset_${name}('
			text += 'value ${field_type}'
			text += ')\n'
			text += '\tclear_' + name + '()\n' 
		} else {
			rfield_type := '[]$field_type'
			
			text += '\t${name}(index int) ?$field_type\n'
			text += '\t${name}_arr() ?$rfield_type\n'
			text += '\t${name}_size() int\n'
			text += '\tadd_${name}(value ${field_type}) &${field_type}\n'
			text += '\tset_${name}(index int, value ${field_type})\n'
			text += '\tclear_' + name + '()\n'
		}

		text += '\n'
	}

	for _, field in m.map_fields {
		name := field.name
		k := field.key_type
		v := field.value_type
		// field_type := 'map[${g.type_to_type(field.key_type)}]${g.type_to_type(field.value_type)}'
	
		text += '\t${name}(key $k) ?$v\n'
		text += '\tset_${name}(key $k, value $v)\n'
		text += '\tclear_${name}(key $k)\n'

		// TODO additional functions
	}

	// TODO handle oneof blocks and extensions!


	text += '\tserialize_to_array() ?[]byte\n'
	text += '\tparse_from_array(data []byte) bool\n'


	text += '}\n'

	return text
}

fn (g &Gen) gen_message_internal(type_context []string, m &Message) string {
	mut text := ''

	m_name := to_v_internal_struct_name(type_context, m.name)
	m_full_name := type_context.join('') + m.name
	m_interface_name := to_v_interface_name(type_context, m.name)

	// Generate for submessages
	for _, sub in m.messages {
		mut context := type_context
		context << m.name
		text += g.gen_message_internal(context, sub)
	}

	text += '\nstruct $m_name {\n'

	if m.fields.len > 0 {
		text += 'mut:\n\n'
	}

	for _, field in m.fields {
		field_type, _ := g.field_type_to_type(&field, false)
		name := escape_name(field.name)

		if field.label == 'optional' || field.label == 'required' {
			text += '\t${name} ${field_type}\n'
			text += '\thas_${name} bool\n\n'
		} else {
			text += '\t${name} []${field_type}\n'
		}
	}

	for _, field in m.map_fields {
		name := field.name
		k := field.key_type
		v := field.value_type
		// field_type := 'map[${g.type_to_type(field.key_type)}]${g.type_to_type(field.value_type)}'

		text += '\t${name} vproto.Map_${k}_${v}\n\n'


		// TODO additional functions
	}

	text += '}\n'

	// Function for creating a new of that message

	text += 'pub fn new_${m_full_name.to_lower()}() $m_interface_name {\n'
	text += '\treturn $m_name{}'
	text += '\n}\n\n'

	// TODO all of this needs to be significantly cleaned up and refactored
	// Move all of the field generating code into the same place for both interfaces
	// and the internal structs

	for _, field in m.fields {
		field_type, is_field_message := g.field_type_to_type(&field, true)

		name := escape_name(field.name)

		if field.label == 'optional' || field.label == 'required' {
			text += 'fn (o &$m_name) ${name}() ?$field_type {\n'
			text += '\tif o.has_${name} {\n'
			text += '\t\treturn o.$name\n'
			text += '\t}\n'
			text += '\treturn none\n'
			text += '}\n\n'

			text += 'fn (o &$m_name) mutable_${name}() ?&$field_type {\n'
			text += '\tif o.has_${name} {\n'
			text += '\t\treturn &o.$name\n'
			text += '\t}\n'
			text += '\treturn none\n'
			text += '}\n\n'
			
			if is_field_message {
				real_field_type, _ := g.field_type_to_type(&field, false)

				text += 'fn (o mut $m_name) set_${name}(value ${field_type}) {\n'
				text += '\to.${name} = ${real_field_type}(value)\n'
				text += '\to.has_${name} = true \n'
				text += '}\n\n'
			} else {
				text += 'fn (o mut $m_name) set_${name}(value ${field_type}) {\n'
				text += '\to.${name} = value\n'
				text += '\to.has_${name} = true \n'
				text += '}\n\n'
			}


			text += 'fn (o mut $m_name) clear_' + name + '() {\n\to.has_${name} = false\n}\n\n' 
		} else {
			rfield_type := '[]$field_type'
			
			text += 'fn (o &$m_name) ${name}(index int) $field_type {\n'
			text += '\treturn o.${name}[index]\n'
			text += '}\n\n'

			text += 'fn (o &$m_name) ${name}_arr() $rfield_type {\n'
			text += '\treturn o.${name}\n'
			text += '}\n\n'

			text += 'fn (o &$m_name) ${name}_size() int {\n'
			text += '\treturn o.${name}.len\n'
			text += '}\n\n'

			if !is_field_message {
				text += 'fn (o mut $m_name) add_${name}(value ${field_type}) {\n'
				text += '\to.${name} << value\n'
				text += '}\n\n'

				text += 'fn (o mut $m_name) set_${name}(index int, value ${field_type}) {\n'
				text += '\to.${name}[index] = ${}value\n'
				text += '}\n\n'
			} else {
				real_field_type, _ := g.field_type_to_type(&field, false)

				text += 'fn (o mut $m_name) add_${name}() &${field_type} {\n'
				text += '\to.${name} << ${real_field_type}{}\n'
				text += '\treturn &o.${name}[o.${name}.len-1]\n'
				text += '}\n\n'

				text += 'fn (o mut $m_name) set_${name}(index int, value ${field_type}) {\n'
				text += '\to.${name}[index] = ${real_field_type}(value)\n'
				text += '}\n\n'
			}

			text += 'fn (o mut $m_name) clear_' + name + '() {\n'
			text += '\to.${name} = []\n'
			text += '}\n\n'
		}
		text += '\n'
	}

	// TODO oneof, maps and similar


	text += 'fn (o $m_name) serialize_to_array() ?[]byte {\n'
	text += '\treturn none\n'
	text += '}\n'

	text += 'fn (o $m_name) parse_from_array(data []byte) bool {\n'
	text += '\treturn false\n'
	text += '}\n'

	return text
}

pub fn (g &Gen) gen_file_text(f &File) string {
	mut generated_text := g.gen_file_header(&f)

	for _, e in f.enums {
		generated_text += g.gen_enum_definition([], &e)
	}

	for _, m in f.messages {
		generated_text += g.gen_message_definition([], &m)
	}


	generated_text += '////////////////////////////////////////'
	generated_text += '// Internal Definitions'
	generated_text += '///////////////////////////////////////'

	// Then generate the actual structs that back the messages
	for _, m in f.messages {
		generated_text += g.gen_message_internal([], &m)
	}

	return generated_text
}

pub fn new_gen(p &Parser) Gen {
	return Gen{&p.type_table}
}