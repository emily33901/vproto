module compiler

fn to_v_field_name(name string) string {
	return name.to_lower()
}

fn to_v_struct_name(name string) string {
	mut new_name := name[0].str().to_upper() + name[1..]
	new_name = new_name.replace_each(['_', '', '.', ''])

	// Get around the capital letters limitations
	mut was_cap := 0
	for i, c in new_name {
		if c >= `A` && c <= `Z` {
			if was_cap > 1 {
				new_name = new_name[..i] + c.str().to_lower() + new_name[i+1..]
			} else {
				was_cap++
			}
		} else {
			was_cap = 0
		}
	}

	return new_name
}

fn to_v_message_name(context []string, name string) string {
	mut struct_name := ''
	
	for _, part in context {
		struct_name += to_v_struct_name(part)
	}

	struct_name += to_v_struct_name(name)

	// TODO when this limitation is removed also do so here!

	struct_name = struct_name.replace_each(['.', ''])

	return struct_name
}

fn escape_name(name string) string {
	if name in keywords_v {
		return name + '_'
	}

	new_name := name.replace_each(['__', '_'])

	return new_name
}

struct Gen {
	type_table &TypeTable
}

fn (g &Gen) gen_file_header(f &File) string {
	// TODO figure out an appropriate module
	// if the file doesnt have an explicit package set

	return '
// Generated by vproto - Do not modify
module vproto_gen

import vproto
'
}

fn (g &Gen) gen_enum_definition(type_context []string, e &Enum) string {
	e_name := to_v_struct_name(type_context.join('') + e.name)
	mut text := '\nenum ${e_name} {\n'

	for _, field in e.fields {
		text += '\t${to_v_field_name(field.name)} = $field.value.value\n'
	}

	text += '}\n'
	
	// TODO helper functions here 
	// https://developers.google.com/protocol-buffers/docs/reference/cpp-generated#enum

	return text
}

enum type_type {
	message enum_ other
}

fn (g &Gen) type_to_type(t string) (string, type_type) {
	if t in valid_types {
		return valid_types_v[valid_types.index(t)], .other
	}

	if _ := g.type_table.lookup_message([], t) {
		if t[0] == `.` {
			return to_v_message_name([], t[1..]), .message
		}

		return to_v_message_name([], t), .message
	}

	if t[0] == `.` {
		return to_v_struct_name(t[1..]), .enum_
	}

	return to_v_struct_name(t), .enum_
}

fn (g &Gen) field_type_to_type(f &Field) (string, type_type) {
	return g.type_to_type(f.t)
}

fn (g &Gen) gen_message_runtime_info(type_context []string, m &Message) string {
	mut text := '\nconst (\n'

	m_name := to_v_message_name(type_context, m.name)
	m_full_name := (type_context.join('') + m.name).to_lower()

	mut fields_block := ''
	mut name_to_number_map := ''
	mut v_name_to_number_map := ''

	if m.fields.len > 0 {
		fields_block = '\t${m_full_name}_fields = [\n'
		name_to_number_map = '\t${m_full_name}_name_to_number = {\n'
		v_name_to_number_map = '\t${m_full_name}_v_name_to_number = {\n'
	} else {
		fields_block = '\t${m_full_name}_fields = []vproto.RuntimeField\n'
		name_to_number_map = '\t${m_full_name}_name_to_number = map[string]i64\n'
		v_name_to_number_map = '\t${m_full_name}_v_name_to_number = map[string]i64\n'
	}

	// TODO should probably also be a map but we cant rn
	// mut number_to_field_func := '\t${m_full_name}_v_name_to_number = {\n'

	for _, field in m.fields {
		field_type, field_type_type := g.field_type_to_type(&field)
		name := escape_name(field.name)

		enum_field_type := if field_type == 'string' || field_type == 'bool' {
			field_type + '_'
		} else if field_type_type == .message {
			'message'
		} else if field_type_type == .enum_ {
			'enum_'
		} else {
			field.t
		}

		fields_block += '\t\tvproto.RuntimeField{\'$field.t\', \'$field_type\', vproto.FieldType.$enum_field_type, \'$field.name\', \'$name\', $field.number},\n'

		name_to_number_map += '\t\t\'$field.name\': i64($field.number)\n'
		v_name_to_number_map += '\t\t\'$name\': i64($field.number)\n'
	}


	if m.fields.len > 0 {
		fields_block += '\t]\n'
		name_to_number_map += '\t}\n'
		v_name_to_number_map += '\t}\n'
	}

	text += name_to_number_map
	text += v_name_to_number_map
	text += fields_block

	text += '\n)\n'



	return text
}

fn (g &Gen) gen_message_internal(type_context []string, m &Message) string {
	mut text := ''

	m_name := to_v_message_name(type_context, m.name)
	m_full_name := (type_context.join('') + m.name).to_lower()

	// Generate for submessages
	for _, sub in m.messages {
		mut context := type_context
		context << m.name
		text += g.gen_message_internal(context, sub)
	}

	text += g.gen_message_runtime_info(type_context, m)

	text += '\nstruct $m_name {\n'

	if m.fields.len > 0 {
		text += 'mut:\n\n'
	}

	for _, field in m.fields {
		field_type, _ := g.field_type_to_type(&field)
		name := escape_name(field.name)

		if field.label == 'optional' || field.label == 'required' {
			text += '\t${name} ${field_type}\n'
			text += '\thas_${name} bool\n\n'
		} else {
			text += '\t${name} []${field_type}\n'
		}
	}

	for _, field in m.map_fields {
		name := field.name
		k := field.key_type
		v := field.value_type
		// field_type := 'map[${g.type_to_type(field.key_type)}]${g.type_to_type(field.value_type)}'

		text += '\t${name} vproto.Map_${k}_${v}\n\n'


		// TODO additional functions
	}

	text += '}\n'

	// Function for creating a new of that message

	text += 'pub fn new_${m_full_name}() $m_name {\n'
	text += '\treturn $m_name{}'
	text += '\n}\n\n'

	// TODO all of this needs to be significantly cleaned up and refactored
	// Move all of the field generating code into the same place for both interfaces
	// and the internal structs

	for _, field in m.fields {
		field_type, field_type := g.field_type_to_type(&field)

		name := escape_name(field.name)

		if field.label == 'optional' || field.label == 'required' {
			text += 'fn (o &$m_name) ${name}() ?$field_type {\n'
			text += '\tif o.has_${name} {\n'
			text += '\t\treturn o.$name\n'
			text += '\t}\n'
			text += '\treturn none\n'
			text += '}\n\n'

			text += 'fn (o &$m_name) mutable_${name}() ?&$field_type {\n'
			text += '\tif o.has_${name} {\n'
			text += '\t\treturn &o.$name\n'
			text += '\t}\n'
			text += '\treturn none\n'
			text += '}\n\n'
			
			if field_type == .message {
				text += 'fn (o mut $m_name) set_${name}(value ${field_type}) {\n'
				text += '\to.${name} = value\n'
				text += '\to.has_${name} = true \n'
				text += '}\n\n'
			} else {
				text += 'fn (o mut $m_name) set_${name}(value ${field_type}) {\n'
				text += '\to.${name} = value\n'
				text += '\to.has_${name} = true \n'
				text += '}\n\n'
			}


			text += 'fn (o mut $m_name) clear_' + name + '() {\n\to.has_${name} = false\n}\n\n' 
		} else {
			rfield_type := '[]$field_type'
			
			text += 'fn (o &$m_name) ${name}(index int) $field_type {\n'
			text += '\treturn o.${name}[index]\n'
			text += '}\n\n'

			text += 'fn (o &$m_name) ${name}_arr() $rfield_type {\n'
			text += '\treturn o.${name}\n'
			text += '}\n\n'

			text += 'fn (o &$m_name) ${name}_size() int {\n'
			text += '\treturn o.${name}.len\n'
			text += '}\n\n'

			if field_type != .message {
				text += 'fn (o mut $m_name) add_${name}(value ${field_type}) {\n'
				text += '\to.${name} << value\n'
				text += '}\n\n'

				text += 'fn (o mut $m_name) set_${name}(index int, value ${field_type}) {\n'
				text += '\to.${name}[index] = value\n'
				text += '}\n\n'
			} else {
				text += 'fn (o mut $m_name) add_${name}() &${field_type} {\n'
				text += '\to.${name} << ${field_type}{}\n'
				text += '\treturn &o.${name}[o.${name}.len-1]\n'
				text += '}\n\n'

				text += 'fn (o mut $m_name) set_${name}(index int, value ${field_type}) {\n'
				text += '\to.${name}[index] = value\n'
				text += '}\n\n'
			}

			text += 'fn (o mut $m_name) clear_' + name + '() {\n'
			text += '\to.${name} = []\n'
			text += '}\n\n'
		}
		text += '\n'
	}

	// TODO oneof, maps and similar


	text += 'fn (o $m_name) serialize_to_array() ?[]byte {\n'
	text += '\treturn none\n'
	text += '}\n'

	text += 'fn (o $m_name) parse_from_array(data []byte) bool {\n'
	text += '\treturn false\n'
	text += '}\n'

	text += 'fn (o $m_name) field_name_to_number(name string) ?i64 {\n'
	text += '\tif name in ${m_full_name}_name_to_number {\n'
	text += '\t\treturn ${m_full_name}_name_to_number[name]\n'
	text += '\t}\n'
	text += '\treturn none\n'
	text += '}\n'

	text += 'fn (o $m_name) field_v_name_to_number(name string) ?i64 {\n'
	text += '\tif name in ${m_full_name}_v_name_to_number {\n'
	text += '\t\treturn ${m_full_name}_v_name_to_number[name]\n'
	text += '\t}\n'
	text += '\treturn none\n'
	text += '}\n'

	text += 'fn (o $m_name) field_from_number(num i64) ?vproto.RuntimeField {\n'
	text += '\tfor i, x in ${m_full_name}_fields {\n'
	text += '\t\tif x.number == num {\n'
	text += '\t\t\treturn ${m_full_name}_fields[i]\n'
	text += '\t\t}\n'
	text += '\t}\n'
	text += '\treturn none\n'
	text += '}\n'

	return text
}

pub fn (g &Gen) gen_file_text(f &File) string {
	mut generated_text := g.gen_file_header(&f)

	for _, e in f.enums {
		generated_text += g.gen_enum_definition([], &e)
	}

	// Then generate the actual structs that back the messages
	for _, m in f.messages {
		generated_text += g.gen_message_internal([], &m)
	}

	return generated_text
}

pub fn new_gen(p &Parser) Gen {
	return Gen{&p.type_table}
}