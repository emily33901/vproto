module vproto