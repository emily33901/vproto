module vproto
